library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
   constant ZERO          : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"03630303230367138303836303b7139323932337b72323232313033763ef1317",
INIT_01 => X"6f330303036f13238337ef0323339303ef2323930303e3032303233333330303",
INIT_02 => X"830383ef036383132323232313676f63672393832383631313672337e31303b7",
INIT_03 => X"6313831363930313631313930323131363138323036f1303ef23036313671313",
INIT_04 => X"936f136f0303ef232303833313e3131363b313239363139383e3136313631363",
INIT_05 => X"63638313b76303936f13ef9303836f1363136f93136fe3939313031313331333",
INIT_06 => X"0303ef23239303e31313836f9313836f13130303ef2323036f1303ef230383e3",
INIT_07 => X"03830333838303ef23131393830383ef232323232323132313939337931313b3",
INIT_08 => X"b303b3676313670337e31303b7671303376f930303ef232303836fe393030323",
INIT_09 => X"139313136313836313839313639313138393232323136fa313676313336f2313",
INIT_0A => X"03833363230363e313933383038303ef23232323139313631363131383231393",
INIT_0B => X"9367138303831323636f136363036393ef23931313232323136f13e313671383",
INIT_0C => X"671313830383630313232323232313671383ef23232323231313932323136fa3",
INIT_0D => X"9393231303b313ef1337e3931303ef13639303ef13372383b313ef931337b303",
INIT_0E => X"936f13636313631393136f9313336393676313136f136f13ef13e3139303ef63",
INIT_0F => X"3767231303b723938323938337232393376f136f13671363e393933333636f93",
INIT_10 => X"ef133723b7ef3723232313931337b7676713371383ef2337b713133763133783",
INIT_11 => X"ef1337e393639363936393e39303ef23efef1337ef1337ef1337ef1337ef1337",
INIT_12 => X"37ef13376fb737ef13376703339313b7e393136fe713ef133793ef139313ef13",
INIT_13 => X"83ef630383ef2323133723339313efef1393379313ef139313ef13ef13376fb7",
INIT_14 => X"1303e31313efef13376fef133763036f932313e3136f938303ef231323631313",
INIT_15 => X"13ef13ef13376f133783e3138303ef13639303ef231323b3b703339323b71323",
INIT_16 => X"13ef133723ef139313ef13ef13376fef139303ef139313ef13ef133723ef1393",
INIT_17 => X"83ef131393ef13ef13376fef1313930383ef139313ef13ef133723ef139313ef",
INIT_18 => X"3cefefef23136f2303ef139313ef13ef133723ef139313ef13ef13376fef1337",
INIT_19 => X"200a4d2020506373200a0a2d64742020520a30204a202025780a00633834304c",
INIT_1A => X"65200a726577642072200a6c2f7568200a4f45657270200a0062200a79696175",
INIT_1B => X"0079252d3f506f740a00640a740a0a787861612020740a7820720a656c4d0a64",
INIT_1C => X"58d874747474747474747474744870e8741c0065640a0a250065650a2928670a",
INIT_1D => X"000000000000000000000000000000000000000000000000000000001074b474",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"277a272524a780012424206c2745068428062064842a2c262e01274700000101",
INIT_01 => X"f007232527f00628266700252a05052700202205272574272627280707072325",
INIT_02 => X"242420f025924584202a2e2c0180f0848020862680260e85078020471c77a706",
INIT_03 => X"8205450414054507f8770705472204078c07262247f00426f022258e07800105",
INIT_04 => X"16f004f02326f02224254507070e07034e04030205940605249605820580056c",
INIT_05 => X"1284458616162604f086f0042545f0058405f00507f0fcf20205430407071787",
INIT_06 => X"2327f024260525d6060324f0050624f007062726f0242625f00727f02425255c",
INIT_07 => X"23254505232227002a8503042523230026282a2c2e2085240302061505060704",
INIT_08 => X"06c3868014078025470c77a70680752507f0842326f024262525f0fa82262780",
INIT_09 => X"050206049607459c074506049606040745842e2a2c01f00f0780140706f08007",
INIT_0A => X"24200584a02786940303052626222700222426280505876687f8870445200303",
INIT_0B => X"84800124242005809000059858270e06f02004070426222401f0876a87800124",
INIT_0C => X"8001052424206e27042220262a2801800120f020202e2c260506052a2801f08f",
INIT_0D => X"f6062406c58607f0051514060727f005180627f0051724c58607f08505170427",
INIT_0E => X"950005d60a05f8050607f0d5170584f680940507f005f004f0051a070627f064",
INIT_0F => X"0780a067a74620f62620e6264720280647f006f00680050496d5d6650766f096",
INIT_10 => X"f005172004f004222e200585011515800001070520f02405050601269a077726",
INIT_11 => X"f00515120600060206ce06c20627f022f0f00515f00515f00515f00515f00515",
INIT_12 => X"04f00515f00404f00515002707861716ec0607f08005f0051504f0050506f005",
INIT_13 => X"26f00c2726f0202207d700060607f0f00505150404f0050506f005f00515f004",
INIT_14 => X"5727100775f0f00515f0f005151a27000520871807f0862627f02005221ef607",
INIT_15 => X"06f005f0051500051525da072627f005987627f02405a0860526061680060722",
INIT_16 => X"05f0051524f0050506f005f00515f0f0050527f0050506f005f0051522f00505",
INIT_17 => X"45f0050605f005f00515f0f00586752726f0050506f005f0051522f0050506f0",
INIT_18 => X"4ef0f0f02401f00027f0050506f005f0051522f0050506f005f00515f0f00515",
INIT_19 => X"555b0053654d7465655b0020656c625349483239617c0030202500643935313e",
INIT_1A => X"637353642072207765775b6c206d65665b4d45786172205b006f425b006e6470",
INIT_1B => X"0074642d0a5220657700616e0a62002e25747262666977292865616465205300",
INIT_1C => X"090b08080808080808080808080b090a0809007820770030007820623a68746c",
INIT_1D => X"000000000000000000000000000000000000000000000000000000000c080908",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"81e5c181e105004181c101d741027404010511007d0191e181c107020010c100",
INIT_01 => X"5f6701c1811f77a141000001a1e5840100e1d1844101e601e181e1a7976701c1",
INIT_02 => X"4181c1df01050405a19111810100df0500d71607b60707050500a70307270603",
INIT_03 => X"a5300414b5c004f0e5f7079004e11400e60041e114df14411fc101e550000100",
INIT_04 => X"275f241f41819f61c101072743e3f0f3906710b10004460006a580a540a530b5",
INIT_05 => X"070506c6000606469f049f4601065f80a5501f9000df55f203140405076717e6",
INIT_06 => X"c1819fe161d001040346069fa046065ff716c1811fc1e1015ff781dfe10141e0",
INIT_07 => X"410105a7c1c18140610313050141c1c091b161e151c104d100414500a003f790",
INIT_08 => X"e506e500e60000070307170603001507035ff481c15f61c101415fb3120181a2",
INIT_09 => X"00940024e58014e500041015e50005d00505119181011fb71700c705c55f6617",
INIT_0A => X"81c1a006e40104829090e50141c18100c1e151d1060595e3f5e3051404819090",
INIT_0B => X"1400014181c10404e40000840501d5a01fe105f505119181011f95e3f5000141",
INIT_0C => X"008100c10141e44100b1a1911181810041c19fc1f1e1d111000105c1b1c15fa4",
INIT_0D => X"f605e1e006e4009f8500d7001781df00d770819f0700e106e4005f0487008701",
INIT_0E => X"1540000505f5e51010055f1517e50615000500059fe0df045fc0d7170081dfd6",
INIT_0F => X"0000e6070600d77607d746070107d720031f109f00000706061516d5b7b71f16",
INIT_10 => X"df870001001f0011918185c58100000007c10000811f110000064100e6170007",
INIT_11 => X"df4500d720d750d700e610e670419fa11f1f4500dfc5009f05005f05001f8500",
INIT_12 => X"001f45009f00009f45000707d7862700e650e75f04005f8500055fc100009fc1",
INIT_13 => X"015f0541015fd1e10703e6d400059f9f45040005051fc100005fc19f45001f00",
INIT_14 => X"2701e590f55f5fc500df5f05000701c007e11607f79f1601418fd1a0a106f605",
INIT_15 => X"005fc19f450040050001e6174181cf3006f7810fe150c6b60006d427068000e1",
INIT_16 => X"c11f0500a11fc100005fc19f45001f5f0705419fc10000dfc11f0500a11fc100",
INIT_17 => X"051fc100005fc19f45001fdf0706f581411fc100005fc19f0500a19fc10000df",
INIT_18 => X"55df9fdf11411fa7411fc100005fc19f8500a19fc10000dfc11f45009f1f0500",
INIT_19 => X"5d7500527820206c5d730025726f6f6f534632206e0000320030006561363200",
INIT_1A => X"7465500a77692f6f615d72006670785d640050746d6f5d50006f5d620061206c",
INIT_1B => X"0065203e004f45207200746f006f002e302079696f6e613a6873640063735200",
INIT_1C => X"0000000000000000000000000000000000000029286f00380029287900656865",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"00060000000000020101020001e11a84000002000100000000fd00e10046ff50",
INIT_01 => X"f900010000f61a0000006e0100001a006f00001a0101fa010000004000000100",
INIT_02 => X"030303fa0002000000020202fc00fb000000000000000000000000e1fe0040e1",
INIT_03 => X"0e070000000600ff0c0ffd00000000020a03000000fb0000f800000002000400",
INIT_04 => X"00f500fd0000eb000000000002f4ffff1c4000020316000100f80514060c060a",
INIT_05 => X"020000c700000000ec00e4000000f5070807fe0000f3fc0ffd000000fd000000",
INIT_06 => X"0000da00000200fe000000ed000000fbff000000df000000feff00e0000000fc",
INIT_07 => X"010100000001003d000000000101003e00000000000200000002c8000000ff40",
INIT_08 => X"0000000000000000e1fe0040e1000040e1e0ff0000cf00000000e2f800020100",
INIT_09 => X"000001000007000003000000000000020000000000fefffe0000000000fe0000",
INIT_0A => X"01014000000000fa010000010000001f000000000000fc06fb00fd0000000100",
INIT_0B => X"00000100000000000201000000000000e900000400000000fff9fafcf9000201",
INIT_0C => X"0001000001010000000000000000fe000200b100020000000001000000fdfbfe",
INIT_0D => X"0ffe0005000000f2ca00fc010000a302000000f5ca0000000000f700c9000000",
INIT_0E => X"0002000002ff00020000fe000000000000000000fd02f3019e07fc0001009f02",
INIT_0F => X"3300001500e100ff00000000e100001be1fa00fa00000000fe0000004000fe00",
INIT_10 => X"d8cd000040da40060406cbcaf90000000000400000c4004033f0ff0002bbb50e",
INIT_11 => X"d0d900f8040a0516050406fa0700b800b9d5d500d5d300d6d200d7d100d8cf00",
INIT_12 => X"30c9d800f04040cad700000000e30000f201f9f40000cedc0000b9000001c900",
INIT_13 => X"00a5020000a50000090000000000a8c4da00000000b0000001c000c7d900ef30",
INIT_14 => X"4000e005fd9ebadd00e1bbdd00000009000000fafffa000000ee000300003f00",
INIT_15 => X"01aa00b1d90012df0000fa000000e302000f00d6000000003b000000003b0000",
INIT_16 => X"00a9e0000094000001a400abd900d3b000000097000001a700afe000009a0000",
INIT_17 => X"008b0001009b00a2d900ca8b00000f00008f0000019f00a6e1000091000001a1",
INIT_18 => X"4cbcb8b400ffc100008500000195009ce200008700000197009fd900c6a0e200",
INIT_19 => X"202c0041742f5365202c007320616f43432d0032200000780038006662373300",
INIT_1A => X"656c4d006f74207264202c00692064202c005220206720200074202c0072626f",
INIT_1B => X"00736220004d457469006120006f002e3830206e726769006573640074654100",
INIT_1C => X"000000000000000000000000000000000000003a68720078003a68740078206e",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
