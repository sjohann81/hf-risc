library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
   constant ZERO          : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"03830383038363831393372393239323232323b723233723231383b763ef1317",
INIT_01 => X"03836f23ef93032333ef930303e383238323b3b3b38303836383032383671383",
INIT_02 => X"2323232323232393b72313676f1363672313032303636723b7e39383376fb383",
INIT_03 => X"6f13ef1363936713138303830383038303830383ef9313638323931393232323",
INIT_04 => X"8313639383e3939313831313331333936f136f93136393931393831313639303",
INIT_05 => X"ef136f936363638393b7631383e393639363936f93ef131383e3936393636393",
INIT_06 => X"93036f1393036fef1383b393e393136333932393639313036f13ef13936f1393",
INIT_07 => X"b76f13ef13936fe31393ef2393138333939383ef139393931313ef331393e393",
INIT_08 => X"2323232323136fa393676393336f23933383336763936703b7e3938337671303",
INIT_09 => X"1363931363938313939313131313639303639303931363931313930323232323",
INIT_0A => X"2323232323136f13671383038303830383038333632363630333ef2313939363",
INIT_0B => X"2323231313932323136fa393671383038303831323636f13636363ef93931313",
INIT_0C => X"8363b39337939337b7131313232323232323232323232313671383ef23232323",
INIT_0D => X"9303b393ef13e393ef1363ef1383b393ef139367131383038303830383038303",
INIT_0E => X"13936363936363936313936f9313b36313671363936f136f13ef13e3ef936393",
INIT_0F => X"03b76723938337231303231303b7232313b76f136f136f9313b333636f139367",
INIT_10 => X"232323232323232323232313931337b7676713371383ef2337b71313376393b7",
INIT_11 => X"93ef93efef1337ef1337ef13ef13ef13ef13b7ef13b7ef13b737b7371337efb7",
INIT_12 => X"13ef133793ef139313ef13ef1337e39363936fef133763e39363936363936363",
INIT_13 => X"63936fef133783ef131393ef13ef1337e39363936363936fef1393ef139313ef",
INIT_14 => X"ef13376f37b7ef13376f23ef139313ef13ef133793ef139313ef13ef1337e393",
INIT_15 => X"13631393ef63ef1323b3b71313efef1393371393ef139313ef13ef13376f37b7",
INIT_16 => X"9393e39313efef13376fe713ef133713ef139313ef13ef13376f13e3136f13ef",
INIT_17 => X"133793ef139313ef13ef13376f139337e393ef136313ef23133383b32313b737",
INIT_18 => X"202025780aefefef23136fef131393ef139313ef13ef133713ef139313ef13ef",
INIT_19 => X"79696175200a4d2020506373200a0020656c6253494830205300633834304c3c",
INIT_1A => X"65200a726577200a642072200a0066200a7568200a4f45657270200a0062200a",
INIT_1B => X"0079252d3f506f740a00640a740a0a787861612020740a7820720a656c4d0a64",
INIT_1C => X"0000000000000000000000000000000000000065640a0a250065650a2928670a",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"2a2929242420e42704844a2409200a262a2c2e84262264222401a74700000101",
INIT_01 => X"2727f024000525260500052925fc272227248787872627277e2727202780012a",
INIT_02 => X"2022242626282e871a2a0180f085868020072700270e80a0479cf72707f08726",
INIT_03 => X"f00bf0858a078001052c2c2b2b2a2a2929242420f005859445260b8b0922242c",
INIT_04 => X"470b940746fcf78705460b0404148417f00b000504e2f7870406470a0b08074a",
INIT_05 => X"f085f00b401884c584179689a4980680068806f00bf08584c590068806e68a06",
INIT_06 => X"84a9f00c8ba9f0f085c5870786840444040408071a8b0ca9f004f08505f00484",
INIT_07 => X"07f004f08505f0f4098c0080840546850a0527000505040c0c04f0098505568b",
INIT_08 => X"2a2e24262c01f08f8780940706f0008707468780140780a5478cf727078075a5",
INIT_09 => X"87f88487fe8447090a0b050b06041607471c0747090416098a0407472e202228",
INIT_0A => X"2e26282a2c01f00480012b2b2a2a2929242420058420041026050026050584e2",
INIT_0B => X"28262e050605242201f08f8480012929242420058094000598580cf009040904",
INIT_0C => X"20ee070c1c090b1b1a048a092226222426282a2c2e202401800120f0262e2c2a",
INIT_0D => X"07c50704f0059084f00596f005c50704f085058001052c2c2b2b2a2a29292424",
INIT_0E => X"8507041007de8887f80707f0d5158704f780859607f005f004f00592f084e0f7",
INIT_0F => X"a7078020e72747a077a7a067a747a0a80747f006f006f0d557e70566f0179580",
INIT_10 => X"2a2c2e262e202224282a2c0585011515800001030520f02605050601261a8777",
INIT_11 => X"07f00bf0f00515f00515f005f085f005f08517f08517f085171b1a1a0409f004",
INIT_12 => X"05f005150bf0050506f005f005159c078407f0f005151c9e078207c48007c08a",
INIT_13 => X"8e07f0f0051545f0050605f005f0051590078e07c68a07f0f08505f0050506f0",
INIT_14 => X"f00515f00904f00515f080f0050506f005f005150bf0050506f005f005159c07",
INIT_15 => X"05960c77f002f08c8087db040cf0f00585150904f0050506f005f00515f00904",
INIT_16 => X"095b140775f0f00515f00005f0051509f0050506f005f0051500041a0cf004f0",
INIT_17 => X"05150bf0050506f005f00515f0050515d689f00516f7f0200507a68600970c0c",
INIT_18 => X"7c00302025f0f0f02601f0f0850675f0050506f005f005150cf0050506f005f0",
INIT_19 => X"006e6470555b0053654d7465655b0025726f6f6f534631316500643935313e4e",
INIT_1A => X"637353642072205b007765205b0069205b6d65205b4d45786172205b006f425b",
INIT_1B => X"0074642d0a5220657700616e0a62002e25747262666977292865616465205300",
INIT_1C => X"000000000000000000000000000000000000007820770030007820623a68746c",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"81c1014181c137c184040201052174115141317d019100f1810107020010c100",
INIT_01 => X"4101dfa1400481a1250004c181fa81f101f1e797d7814101f74101f10a000141",
INIT_02 => X"219181117161318a005101001f050500e51705b7050500a70307270703dfd781",
INIT_03 => X"1f1b5f09f5500001004181c1014181c1014181c1df0009050bf1060505918141",
INIT_04 => X"0b1bf6c00bf5f7061b0b0504d41487249f2b409000f6f707f0900b001bfa001b",
INIT_05 => X"df095f09800405040700044b0bd730d780d7509f041f094b0bd730d780f6d740",
INIT_06 => X"4b0b9fa04b0b5f9f0907970184f4f0809410f100094b000b1ff45f090a9ff414",
INIT_07 => X"039ff49f090a9f8a051c40dc140905a7090cc100090c0001a0f45f2009d00904",
INIT_08 => X"9111413181011fb71700c705c55fd717f507f500f60000070307170703001507",
INIT_09 => X"f7ea97f79b07f914909000940024f78014f700041015f7000505d00571615121",
INIT_0A => X"113121918101df090001c1014181c1014181c1a0098a0a2bc19580c1060597ea",
INIT_0B => X"e1d111004105c1b1019fa4140001c1014181c10404240000840535dfa005f505",
INIT_0C => X"c14724e000007000000505059111918171615141312181010001c15fc11101f1",
INIT_0D => X"050794001fcc34141f0074df4b0794001fca040001004181c1014181c1014181",
INIT_0E => X"07050607000507f7a510101f1515a70715000705001fe05f045fc0341f14fcf7",
INIT_0F => X"070000f7070700e77707e747070107e720031f109f00df1517e7b5b51f171500",
INIT_10 => X"918171311161514121918185c50100000003010000c15f110000060100f71700",
INIT_11 => X"505f05df1f0500dfc5009fcb1fca9f0a1f0700df87009f870000000000009f00",
INIT_12 => X"015f0500051f0100001f01df4500fb40fb209fdf050004fb00fb2077fb5077fb",
INIT_13 => X"fb509fdf0500059f0100009f015f4500fb20fb6077fb30df5f0b059f0100009f",
INIT_14 => X"1f4500df00009f45005fab9f0100009f015f8500051f0100001f01df4500fb70",
INIT_15 => X"300705f41f059f0b87840300055f9f4504000505df010000df019f45005f0000",
INIT_16 => X"0024f590f55f9fc5005f09001f850005df010000df019f450080140cfc1f14cf",
INIT_17 => X"0500059f0100009f015f45005f0504003b198f3007f9cfd7509706e40c290080",
INIT_18 => X"00003200309f5f9f11019fcf0b0cf59f0100009f015f0500051f0100001f01df",
INIT_19 => X"0061206c5d7500527820206c5d73007320616f43432d39207000656136320055",
INIT_1A => X"7465500a77695d77006f615d72006c5d6670785d640050746d6f5d50006f5d62",
INIT_1B => X"0065203e004f45207200746f006f002e302079696f6e613a6873640063735200",
INIT_1C => X"0000000000000000000000000000000000000029286f00380029287900656865",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"01010202020203001a84e10000031a02010101010002000002fd00e10045ff50",
INIT_01 => X"0000f6006c000000016d000000f8000000004000000000000400000000000301",
INIT_02 => X"05040404030303c80003fb00fc0000000000000000000000e1fe0040e1fa0000",
INIT_03 => X"fa00f30000020005000202020303030304040404f70000040000000000030303",
INIT_04 => X"0000000600fc0ffd000000fd00000000fd00020000040ffdff00000200020300",
INIT_05 => X"e200f00002000000c800000000f20706070a07f400e8000000f6060805020e06",
INIT_06 => X"0000fb000000fedc00000001eaffff0a4000000306000100fdffe10000fdff00",
INIT_07 => X"e1f4ffd30000f5fd00003d0000000000000000400000000100ffd9410002fe00",
INIT_08 => X"0202030302fcfffe0000000000fe00000000000000000000e1fe0040e1000040",
INIT_09 => X"f900fcfb00fdff00010000000100000700000300000000000000020001030303",
INIT_0A => X"0001010000fef70000040102020202030303034000000005000021000000fa02",
INIT_0B => X"0202000002000202fcfbfe00000200010101010000030100000001e700000400",
INIT_0C => X"0203410500010000000000000202010101010101010302fd000401b400030302",
INIT_0D => X"fe000000efc7ff00a30201f0c7000000f2c60000030000000001010101020202",
INIT_0E => X"00000002000000ff000002fe000000000000000000fe02f5019f07ffa000020f",
INIT_0F => X"0e3300001500e100ff00000000e100001be1fa00fa00fc0000004000fd000000",
INIT_10 => X"0505050706070707070606cac9f80000000001400000c0004033f0ff0002bbb5",
INIT_11 => X"06b100b1cfd600cfd400d0d3d1d2d1d1d2d000d2ce00d3cc000000000040d540",
INIT_12 => X"00c6e00000b0000001c100c8d900f4062006f6cadd0022f60520040318050b16",
INIT_13 => X"0a07eabee20000a8000100b900c1d900ee072006050a07efc80000ad000001be",
INIT_14 => X"b6d800e24040b7d700e400a1000001b200bae20000a4000001b500bcd900e807",
INIT_15 => X"0200003f92029109010000000094b1da000000009b000001ac00b4d900e13030",
INIT_16 => X"0040d205fd8aa7dd00d40000a9dc000092000001a300abd9000a00fcfffd00e0",
INIT_17 => X"e00000870000019800a0d900e2df0000fd00d502000fc6000001000000003b3b",
INIT_18 => X"0000780038bdb9b500ffc4ff00000f8200000193009be100008500000196009d",
INIT_19 => X"0072626f202c0041742f5365202c000a2d64742020520032200066623733004c",
INIT_1A => X"656c4d006f7420200072642020006c202000642020005220206720200074202c",
INIT_1B => X"00736220004d457469006120006f002e3830206e726769006573640074654100",
INIT_1C => X"000000000000000000000000000000000000003a68720078003a68740078206e",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
