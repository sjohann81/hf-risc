library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
   constant ZERO          : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"3c00afafafafafaf3caf8c273c27038cac8f3c30240caf273c000010000c273c",
INIT_01 => X"1400008f8faf008e001000008f00102c008faf008faf000000008f8f8f2608af",
INIT_02 => X"001400008faf240c8faf00000c8f248f00142c008faf008faf0000008f8f8f00",
INIT_03 => X"2c272400038c3c1030008c3c30038c3c0003ac3c1030008c3c27038f8f8f8f8f",
INIT_04 => X"2406a01626900202000c0200020c020200260800003c001000afafafafafafaf",
INIT_05 => X"10300010a20826a00827038f8f8f8f8f8f028fa014a000242480800210a00224",
INIT_06 => X"1400000000140000001000142400000004001000082404241000000300140000",
INIT_07 => X"0c003a24040027038f00008f00000c0004af04af272408000800030003001400",
INIT_08 => X"2602000c0024240824240000afafafafafafaf272408000827038f00008f0000",
INIT_09 => X"27038f8f8f8f8f8f028f0008001024142c24142c24142e24100010000c00102a",
INIT_0A => X"8f8f00140080002732260c00100083240cafaf27270008260c24240c240c0012",
INIT_0B => X"08240c27038f8f00140080002732260c00100083240c27020014afaf2c272703",
INIT_0C => X"048c0010ac000024000030000000008c8cac34008cac002408243c0024000002",
INIT_0D => X"ae348f8e000c000c00000c0000240cae30afaf00248e3caf2700030008ac3400",
INIT_0E => X"0226322612000c00000c0000000c3024ac30afafafaf0027248c3c2703308f8f",
INIT_0F => X"8e000c24ae30afafaf0024af8e3caf272703ac8f8f8f348f8c3c001626a2000c",
INIT_10 => X"270824ac348f8f8f8f8f8c3c16260c82000c00000c0000260cae00008eae3424",
INIT_11 => X"00102402003c02000c24020c002400000c24000cac00248cacafafaf34278c3c",
INIT_12 => X"27033c008f8f8f300c3c24000002000c24020c002400000c24240c27038f8f8f",
INIT_13 => X"140082260c26243c00140082260c24000c260cafafafafafafafafaf3caf3427",
INIT_14 => X"82260c26243c00140082260c26243c00140082260c26243c2424242700240c00",
INIT_15 => X"240c00140082260c26243c00140082260c26243c00140082260c26243c001400",
INIT_16 => X"82260c2624003c0c00140082260c26243c0000008c0024003c102c26000c000c",
INIT_17 => X"0c2610000c24123608a03c02000c00140082260c26243c3c3c08ae000c001400",
INIT_18 => X"24003c0c00140082260c26243c00083c0c00140082260c26243c260824103226",
INIT_19 => X"0c90022400140082260c2426020c3c240c020026002418000c00140082260c26",
INIT_1A => X"18000c00140082260c26243c2608240c0016240c000c90022600120012240c00",
INIT_1B => X"300c022626120012240c24000c300c023200140082260c2426020c3c240caf00",
INIT_1C => X"0c00140082260c2624003c0c00140082260c26243c260826240c0016240c000c",
INIT_1D => X"0c00140082260c26243c24083c1424a00202301a000c00140082260c2624003c",
INIT_1E => X"24263c0c0200140082260c263c241224083c0200140082260c26243c3c00083c",
INIT_1F => X"00162402a0269000123c000027a3a3a3a3a3a324a300000024a324140082260c",
INIT_20 => X"26243c02088f260caf27082712270c33162402a02690021227273c0012270c00",
INIT_21 => X"140082260c26243c3c080016240c0016260c2400142c2400922600140082260c",
INIT_22 => X"08a0083c088f001402260c2416320c002624102c24020c2412320c2632082600",
INIT_23 => X"62666a6e72767a6c283c0800140082260c24263c0c022600140082260c263ca0",
INIT_24 => X"200a2062200a79696175200a3031442d647420520a7874706c68643935313337",
INIT_25 => X"2d2e612020740a7820720a746577200a00666d200a00646d200a4d456d2f7270",
INIT_26 => X"0000000000000000000065610a0065650a20202928670a206d670a740a652000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000001000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"1180b3bfa0b0b1a212b242bd02bde06262bf03428400bfbd048000000000bd1d",
INIT_01 => X"404300a3a2a2002200405000a200404200a2a200a2a244526200a2a4a35200a0",
INIT_02 => X"00405000a2a20500a4a2530000b305a400404200a2a200a2a2446200a3a4a200",
INIT_03 => X"42bdc200e04202404200620342e0420200e044024042006203bde0b0b1b2b3bf",
INIT_04 => X"022082008462a222400040404000200080b500a08015a040c0b0b1b4b5bfb2b3",
INIT_05 => X"60a300a0820084a000bde0b0b1b2b3b4b560bf85406683846386656040806383",
INIT_06 => X"6003438500e08500006003e042a40500a00040050002a00340a400e004a04405",
INIT_07 => X"00051010a104bde0b05062bf10000000a0b080bfbd0300000080e000e000c005",
INIT_08 => X"523010004051150014130000b1bfb0b2b3b4b5bd06000000bde0b05062bf1000",
INIT_09 => X"bde0b0b1b2b3b4b500bf40004055516063436063436023515400530000004042",
INIT_0A => X"b0bf0080004470a3101000008000a40600bfb0a5bd1000520004040004000040",
INIT_0B => X"000400bde0b0bf0080004470a3101000008000a40600a5008040bfb082bdbde0",
INIT_0C => X"816500e0664504e704c8a502020405666565a5026565a9080009030007040400",
INIT_0D => X"0363bf0300000400110400041104000291b1bf43030210b0bd00e0000065a500",
INIT_0E => X"113131312004001204000412a000d1046292b0b1b2bf47bd076203bde042b0b1",
INIT_0F => X"23a000042392b0b2bf7313b32311b1bdbde062b0b1b242bf6203001110020000",
INIT_10 => X"bd00046242b0b1b2b3bf62031110000404001204000412110022531222236304",
INIT_11 => X"00436302110302400004220011040240000400004365054343b0b1bf63bd4302",
INIT_12 => X"bd201900b0b1bfc600050446110240000422001104024000040400bde0b0b1bf",
INIT_13 => X"80000410001004100080000410000400001000b1b2b3b4b5b6b7bebf10b004bd",
INIT_14 => X"041000100410008000041000100410008000041000100410161217b100040000",
INIT_15 => X"0400008000041000100410008000041000100410008000041000100410008000",
INIT_16 => X"0410001004401000008000041000100410004000426263020360430240000000",
INIT_17 => X"0010400000040010006210740000008000041000100410131000620000008000",
INIT_18 => X"0440130000800004100010041040001000008000041000100410940004608310",
INIT_19 => X"0044701300800064730004730000130400a20215024240000000800064730073",
INIT_1A => X"4000000080000410001004107300040000770400000044707300720077040000",
INIT_1B => X"840015b5949200b614000440008400157000800004100004106000100400b440",
INIT_1C => X"0000800064730073044013000080000410001004109400b5040000b604004000",
INIT_1D => X"0000800004100010041004001055424300b043a0000000800064730073044013",
INIT_1E => X"0410100080008000041000101004800400106000800004100010041013400010",
INIT_1F => X"002242144310639060041400a2b4a3a5a0a2a405a514141405a5058000041000",
INIT_20 => X"7304137400a29400a2a200de60a500c4224214431063b060a2de150060a50000",
INIT_21 => X"8000a4b500b50415100000b00400001310000400404282000413008000647300",
INIT_22 => X"0040001000b400407e730004b01000401004606343000004b0100010b5001500",
INIT_23 => X"6165696d717579296e1000008000041000041010008094008000041000101040",
INIT_24 => X"445b006f425b006e6470555b31376520656c6249487975716d69656136323236",
INIT_25 => X"2d2e726266697729286561612072205b006965205b007565205b005070206172",
INIT_26 => X"00000000000000000000782064007820627c203a68746c006972700a62736200",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"f080000000000000010000fff00000000000f0ff780100ff012800ff0002ff50",
INIT_01 => X"ff10000000000000000010000000006100000000000010101000000000780000",
INIT_02 => X"00ff100000006101000010000100610000ff6100000000000010100000000000",
INIT_03 => X"00ffff000000f0ff000000f0000000f0000000f0ff000000f000000000000000",
INIT_04 => X"0000ffff000018108000282028002088a01100a0880098009000000000000000",
INIT_05 => X"00001000000000000000000000000000001000ffff001000ff000020000010ff",
INIT_06 => X"ff18102000003810100018ffff38280000000028000000000010000020ff1028",
INIT_07 => X"00280000ff200000001010001830008000000000ff0000100010000000000028",
INIT_08 => X"0080810020ff00010000908000000000000000ff000030000000001010001830",
INIT_09 => X"0000000000000000100020018800ffff00ffff00ffff00ff0000000000000000",
INIT_0A => X"000000ff00001000ff0000800000000000000000ff8101ff0000000000000000",
INIT_0B => X"0100000000000000ff00001000ff000080000000000000208000000000ff0000",
INIT_0C => X"ff000000001026ff263000161620280000000010000028ff01fff01000262620",
INIT_0D => X"00000000200126012626012622000100ff000010ff00f000ff00000001000000",
INIT_0E => X"8800ffff00260126260126228001ff0000ff0000000010ffff00f00000000000",
INIT_0F => X"0080010000ff00000018ff0000f000ff000000000000000000f000ff00002001",
INIT_10 => X"0000000000000000000000f0ff00010026012626012622000100109100000000",
INIT_11 => X"0000001012b18088010080018e001488010020010018ff000000000000ff00f0",
INIT_12 => X"00004020000000ff01400030321088010080018e001488010000010000000000",
INIT_13 => X"ff0000000012000000ff0000000000000212000000000000000000000000e1ff",
INIT_14 => X"00000012000000ff0000000012000000ff0000000012000000000000a0000000",
INIT_15 => X"000000ff0000000012000000ff0000000012000000ff0000000012000000ff00",
INIT_16 => X"000000130098000100ff000000001200000000000010131000ff00ff80000000",
INIT_17 => X"00ffff00000001d002000018a00000ff0000000012000040000200000100ff00",
INIT_18 => X"0080000100ff000000001200009802000100ff00000000120000000200010300",
INIT_19 => X"01ff100000ff0000000000132001000000a8110011ffff000100ff0000000013",
INIT_1A => X"ff980100ff000000001300000003000000ff00000001ff100000000000000000",
INIT_1B => X"ff012000000000000000002001ff0120ffa8ff000000000013200100000000f0",
INIT_1C => X"0100ff00000000130080000100ff00000000120000000300000000ff00002001",
INIT_1D => X"0100ff00000000120000000200ff000010a800fe000100ff000000001300a800",
INIT_1E => X"001300012000ff00000000130000fe000200f800ff0000000013000040980300",
INIT_1F => X"00ff0098000000180040988000000000000000ff001c12260000ffff00000000",
INIT_20 => X"130000180200000000000400fe0001ffff00980000001800000040f0fe000120",
INIT_21 => X"ff00000000130000000200fe000000ff000000000000ff00000000ff00000000",
INIT_22 => X"03000400020000ff10000000ffff00200000ff00ff20010000ff0000ff040000",
INIT_23 => X"3964686c7074780075000200ff0000000000130001200000ff00000000120000",
INIT_24 => X"5d50006f5d620061206c5d7536206300726f6f53467a76726e6a666237333135",
INIT_25 => X"3e0079696f6e613a6873640064695d77006c6d5d66006d6d5d64005220646d6f",
INIT_26 => X"0a0a0a0a0a0a0d0a0e0029286100292879000000656865006e6172006f007900",
INIT_27 => X"0a0a0a0a0e0a0c0a0f0a0a0a0a0a0a0a0a0a0a0a0a0c0a0a0a0a0f0a0a0a0a0a",
INIT_28 => X"000000000000000000000000000000000001000b0a0b0a0a0a0a0a0a0a0a0a0a",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"00253034102428187d2c50c8001808e0f01400ff400814e87d2500ff0060fc00",
INIT_01 => X"e32b00181c1c005000292b0010001ea8001418001c142321210014181c403314",
INIT_02 => X"00d92b001014a80a141021000810a81400e4a8001418001c1423210014181c00",
INIT_03 => X"23d0fe0008e000fc40001000400810000008e000fc80001000380824282c3034",
INIT_04 => X"2d1afff20123212325bc252525eb252525e491252500252e25141824282c1c20",
INIT_05 => X"0201250701a00200ad300814181c202428252cfff9012b01ff00002509002bff",
INIT_06 => X"f942252300032b25250a40f8ff2b400008001940d2201f01102b000840fb2142",
INIT_07 => X"c6230101f5231808102126142325c6250d100c14e801d825e125080008000342",
INIT_08 => X"0121006725c908230d0a2525182c141c202428d001c625c61808102126142325",
INIT_09 => X"300814181c202428252c251c250da9ea1a9fec1abff00ad00e00100074001410",
INIT_0A => X"303400f800002110ff0167250a00100a7d343010c80220ff6708206708670008",
INIT_0B => X"6930673808303400f800002110ff0167250a0010107d10252516343010c83808",
INIT_0C => X"e9900008902503ff002401030040c29080900240909024fd9efb002508030025",
INIT_0D => X"90081c90258103810003810002038190ff181c24f7900014e00008008b900400",
INIT_0E => X"2101ffff0a038100038100022581ff0390ff1014181c24e0f790002008ff1418",
INIT_0F => X"9025810690ff141c2424f720900018d8200890101418081c900000fb01002581",
INIT_10 => X"28130a900814181c20249000fc01810003810003810003408190248090900802",
INIT_11 => X"0006b525006b2525a70325a700020025a70125a79024fd909014181c09e09000",
INIT_12 => X"2008002514181cffc5000825002525a70725a700060025a70504a7200814181c",
INIT_13 => X"fb0000016744440000fb000001670a00202c065c6064686c7074787c00580080",
INIT_14 => X"000167780a0000fb00000167680a0000fb00000167500a0007100850250a6700",
INIT_15 => X"0a6700fb00000167c00a0000fb00000167ac0a0000fb00000167980a0000fb00",
INIT_16 => X"0001674c0a25000c00fb00000167d40a0000080000215c8000c136be25740074",
INIT_17 => X"74fffb00702d6790fb000321257400fb00000167e40a0000008900000c00fb00",
INIT_18 => X"0a25000c00fb00000167d40a0025ea000c00fb00000167d40a0001f42a14ff01",
INIT_19 => X"62ff210100fb0000016720342562000a6721001002ff5e000c00fb0000016724",
INIT_1A => X"28250c00fb00000167240a000148206700f620670062ff210100d7000c206700",
INIT_1B => X"ffa7210101bd000d0167202562ffa721ff25fb0000016720342562000a675025",
INIT_1C => X"0c00fb00000167240a25000c00fb00000167d40a00017d01206700f520672562",
INIT_1D => X"0c00fb00000167d40a000a8a00fd01002521ffdb000c00fb000001673c0a2500",
INIT_1E => X"2004004b2500fb0000016714000ab60a8a000900fb000001670c0a000025c500",
INIT_1F => X"00f8012b0001002167002b2518171513121614b5110202026b10b1fb00000167",
INIT_20 => X"38200021f5540167541008017410f0fff8012b0001002154100100258410f025",
INIT_21 => X"fb00000167382000008900fa7c6700f601672e00025fe000001000fb00000167",
INIT_22 => X"fd000e00895000092a10677cf5ff6725012ef65fe025a77c0dff6701ff491000",
INIT_23 => X"3863676b6f7377006c008900fb000001672004004b250100fb00000167fc0000",
INIT_24 => X"202c0074202c0072626f202c0032200020616f432d0077736f6b676338343034",
INIT_25 => X"20002e6e726769006573640061742020006c2020200070202020004f45752067",
INIT_26 => X"2020202020205020d8003a6874003a687400000078206e00676d6f006f007400",
INIT_27 => X"202020202c204c200c2020202020202020202020201820202020442020202020",
INIT_28 => X"000000000000000000000000000000000300003c20a020202020202020202020",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
