library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
   constant ZERO          : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"af00afafafafafaf3caf8c273c27038cac8f3c30240caf273c000010000c273c",
INIT_01 => X"008faf0000008f8f8f000800008f8f8f001000008f8faf008e001000008f263c",
INIT_02 => X"3c1030008c3c27038f8f8f8f8f0008af240c8faf00000c8f248f00142c008faf",
INIT_03 => X"a008001400afafafafafafafaf2c272400038c3c1030008c3c30038c3c0003ac",
INIT_04 => X"8000100002a226a226242606020802a21226900002000c0200020c022600003c",
INIT_05 => X"00242400030008000000103000100027038f8f8f8f8f8f8f028fa008a0242480",
INIT_06 => X"00af04af00002700030000140008000000001400100000000800000400102410",
INIT_07 => X"2408000827038f8f27088f8f0008000c0000080016000c000000000400082404",
INIT_08 => X"00102c240824102c2400142c2410001000000c2424240000afafafafafafaf27",
INIT_09 => X"038f8f8f8f8f8f028f00142a2602000c000008260c24240c240c001200142408",
INIT_0A => X"2702240c0010afaf2c2727038f8f2708320c261000800027000cafaf24272727",
INIT_0B => X"038f8f0008260c0010008200afaf2727038f8f2708320c26100080002700240c",
INIT_0C => X"243c002400000003ac34008c3c0003ac00248c3c0003ac00008cac34248c3c27",
INIT_0D => X"afaf2700030014ac00240000008c003000008c00ac34008cac00340800048c24",
INIT_0E => X"00240c000caf3030afafaf2727038f328f000c000c000c00000c0000240c300c",
INIT_0F => X"0c000c240c000c30afafaf2727088f8f8f8f2608a2000c001202000c00000c00",
INIT_10 => X"24000caf0cafaf272708248f8f8f000c0016260c8226000c00000c0000240c00",
INIT_11 => X"0002000c24020c002400000c24240c00142402003c02000c24020c002400000c",
INIT_12 => X"3c0caf0cafafafafafafafafaf342727038f8f8f27033c008f8f8f300c3c2400",
INIT_13 => X"0c260c240c3c240c3c240c3c240c3c240c3c240c3c2600260c3c240c3c240c3c",
INIT_14 => X"240c3c00162424102a120008000c240c3c0016241224122424102a1224000c00",
INIT_15 => X"ae000c000c243c000c240c3c001624120008000c000c243c000c000c243c000c",
INIT_16 => X"0c00143200000c2610000c02a0023600003c0c240c3c3c0008000c240c3c3c08",
INIT_17 => X"020c240c3c00123c080002240c3c3c26083c08240c3c020c260c243c16260824",
INIT_18 => X"27a0082600902700021002243c0024a3a3a300a300a300a324a324a324240c3c",
INIT_19 => X"32021424a00027a008260090270202100200261002243c00270c00021424a000",
INIT_1A => X"9002242400260c020c260c001000028faf020c000c243c3c0c240c3c0208270c",
INIT_1B => X"27240c3c0008270c00102c240090032400240c3c021626020c262616020c000c",
INIT_1C => X"706c6864393531333762666a6e72767a6c282408a0003c10002608240c3c0317",
INIT_1D => X"646d200a4f457270200a2062200a79696175200a0a3032532d647420520a7874",
INIT_1E => X"28670a6520206d670a740a2e612020740a7820720a746577200a00666d200a00",
INIT_1F => X"0000000000000000000000000000000000002d0065610a0065650a7c2e202029",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"a080b1bfa0b2b3a210b042bd02bde06262bf03428400bfbd048000000000bd1d",
INIT_01 => X"00a2a2446200a3a4a250006200a2a4a300404300a3a2a2006200405200a21013",
INIT_02 => X"024042006203bde0b0b1b2b3bf0000a20500a4a2510000b105a400404200a2a2",
INIT_03 => X"a000c040a0b0b2b3b4b5bfb1b642bdc200e04202404200620342e0420200e044",
INIT_04 => X"6200408320000342500203618000000280504255624000c040c00060b5a08015",
INIT_05 => X"a4020300e0050004440060a300a000bde0b0b1b2b3b4b5b620bf820065846385",
INIT_06 => X"04b081bfa080bd00e06080c0050002628500e08540000002000500a0006063e0",
INIT_07 => X"06000000bde0b0bfbd00b0bf020000004002000000000003400000a1400010a1",
INIT_08 => X"004042920082404282006043425440534000001514130000b2bfb0b1b3b4b5bd",
INIT_09 => X"e0b0b1b2b3b4b500bf0040223150100040100031000404000400002000959200",
INIT_0A => X"a50004008040bfb082bdbde0b0bfa30010001080004470a30000bfb006a5bdbd",
INIT_0B => X"e0b0bf000010000080000480bfb0bdbde0b0bfa30010001080004470a3000600",
INIT_0C => X"09030006040400e0624200620300e0624404620300e0436400434363044302bd",
INIT_0D => X"b0bfbd00e000c06504c6a7040465a2420205620265a5026565a9a50000816507",
INIT_0E => X"120400a000b0d192b1b2bfbdbde0b002bf400000000400100400041004009000",
INIT_0F => X"0011000400a00091b0b1bfbdbd00b0b1b2bf1000020000001111040012040004",
INIT_10 => X"040000b000b1bfbdbd0004b0b1bf000000111000041104001104000411040000",
INIT_11 => X"1102400004020010040240000404000043630211030240000402001004024000",
INIT_12 => X"1200b100b4b5b6b7beb0b2b3bf04bdbde0b0b1bfbd201900b0b1bfc600050446",
INIT_13 => X"0044008400048400048400048400048400048400047300440013840004840004",
INIT_14 => X"8400040022020240222240000000840004002202220222020240222202400000",
INIT_15 => X"2200004000840400008400040022022200000000400084040000400084040000",
INIT_16 => X"00004002400000944000002054b0310040110084000415400000008400040400",
INIT_17 => X"0000840004000004000020840004111000040084000400001000840480100004",
INIT_18 => X"a6c30031e263a7a320c03004050002b0a0a210a210a210a202a202a202840004",
INIT_19 => X"843056426082a4830031e263a7a320803000944030161500a5000030444260c2",
INIT_1A => X"44b1171e00c4002000440000404534a5a280004000840416008400043000a500",
INIT_1B => X"de8400040000de00004042820044d11700840004b1b7b56000b5b5be60000000",
INIT_1C => X"716d696561363232366165696d717579296e630082740480713100840004d1d7",
INIT_1D => X"7565205b4d456172205b006f425b006e6470555b0031326520656c6249487975",
INIT_1E => X"68746c7362006972700a622e726266697729286561612072205b006965205b00",
INIT_1F => X"0000000000000000000000000000000000002d007820640078206200007c203a",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"0090000000000000010000fff00000000000f0ff780000ff012800ff0002ff50",
INIT_01 => X"00000010100000000010001000000000000010000000000000000010000078f0",
INIT_02 => X"f0ff000000f0000000000000000000006100000010000000610000ff61000000",
INIT_03 => X"0000b00088000000000000000000ffff000000f0ff000000f0000000f0000000",
INIT_04 => X"000000102000ff000000ff00980090ff0000001010a00028202800200e909800",
INIT_05 => X"3800000000280020100000000000100000000000000000001000ff000000ff00",
INIT_06 => X"100000001810ff0000101000280010182000003800181010002800000000ff00",
INIT_07 => X"0000300000000000000000001000300020100000003000282080300020000000",
INIT_08 => X"000000ff01ff0000ff000000ff009000200000000000888000000000000000ff",
INIT_09 => X"00000000000000100000ff0000808100908101ff00000000000000000000ff01",
INIT_0A => X"002000008000000000ff000000000001ff00000000001000800000000000ff00",
INIT_0B => X"0000000001000010000000800000ff000000000001ff00000000001000800000",
INIT_0C => X"fff010002626000000000000f000000010ff00f00000001800000000ff00f000",
INIT_0D => X"0000ff000000ff0026ff282620001000102e002e0000100000280001000000ff",
INIT_0E => X"220001800100ffff000000ff000000000080012001260126260126220001ff01",
INIT_0F => X"01890100018001ff000000ff0001000000000001002001000088260126260126",
INIT_10 => X"00200100010000ff000000000000000100ff0001000026012626012622000100",
INIT_11 => X"3210880100800186001480010000010000001012b18088010080018600148001",
INIT_12 => X"00020000000000000000000000e1ff000000000000004020000000ff01400030",
INIT_13 => X"000e010f01000f01000e01000e01000e01000e01000f800e01000e01000e0100",
INIT_14 => X"0f010000ff0000000000880200010f010000ff00000000000000000000880000",
INIT_15 => X"00000188010f0000010f010000ff00001803000188010f000001a0010f000001",
INIT_16 => X"00000003a00000ff000000a00010d080a000000f010040a80200010f01000002",
INIT_17 => X"20010f010000ff000220f80f010040000200020f0100200100010f00ff000200",
INIT_18 => X"000003003000001818003000408800000000120014001600ff000000ff0f0100",
INIT_19 => X"ff20ff00001800000300200000181800201000ff100040a000012030ff000018",
INIT_1A => X"00100000a80f0120010e0100ff101000008801a0010f0000010f010010030001",
INIT_1B => X"000f010000030000000000ff00001000f00f010010ff002001ff000020010001",
INIT_1C => X"726e6a6662373331353964686c70747800750003002000fe2000030f010010ff",
INIT_1D => X"6d6d5d6400506d6f5d70006f5d620061206c5d750036207000726f6f53467a76",
INIT_1E => X"6568650079006e6172006f0079696f6e613a6873640064695d77006c6d5d6600",
INIT_1F => X"0000000000000000000000000000000000003e00292861002928790000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"14212834102c30187d2450c8001808e0f01400ff40fc14e87d2100ff0051fc00",
INIT_01 => X"001c1423210014181c213c210014181c00082b00181c1c0050002d2b00104000",
INIT_02 => X"00fc80001000380824282c3034002214a8fe14102100fc10a81400dda8001418",
INIT_03 => X"00a621032110181c20242c142823d0fe0008e000fc40001000400810000008e0",
INIT_04 => X"0000082b2100ff01022dff05218421ff040123212321b1212121d92140212100",
INIT_05 => X"2b0121000842b2402100020100082130081014181c202428212cff9c0101ff00",
INIT_06 => X"231006142121e8000821210242cb42252300032b08212140bf4000050006ff09",
INIT_07 => X"01bd21bd1808101418bd101423f821bd2123f8000c21bd232121210f21e8010e",
INIT_08 => X"00031ac9309f031abf00190ad0242126210067080d0a21211c2c1418202428d0",
INIT_09 => X"0814181c202428212c00d7100121005a210234ff5a08205a085a0008000da930",
INIT_0A => X"1021305a2103343010c8380830341049ff5a010500002110217034300a10c830",
INIT_0B => X"0810140075015a21050000211410e8380830341064ff5a010500002110211070",
INIT_0C => X"fb00210803000008900800900000089024f790000008902400909009fd900018",
INIT_0D => X"1014e8000800e79003ff240040902501c203800090024090902404a7000390fd",
INIT_0E => X"02039a218c10ffff14181ce0180810ff142193219a039a00039a0002039aff8c",
INIT_0F => X"8c8093069a218cff14181ce020931014181c01e700219a000621039a00039a00",
INIT_10 => X"0121bd1481181ce020130a14181c009300fc019a0040039a00039a0003029a00",
INIT_11 => X"002521bd0725bd00060021bd0504bd001cb525006b2521bd0325bd00020021bd",
INIT_12 => X"00185c06686c7074785860647c0080200814181c2008002114181cffd4000825",
INIT_13 => X"67ac71187100047100f07100d87100c87100b071006821ac7100a07100887100",
INIT_14 => X"2c710000cf667517716221f200002c710000dd4265623855700f65bf64216700",
INIT_15 => X"0000002171a40000002c710000b8771821870000217194000000217174000000",
INIT_16 => X"5a0011ff210067ff0b006321002190212103673c71000021ca00002c7100006c",
INIT_17 => X"21415c71000071006c21095471000001d2006c6c710021410171b400f101d22a",
INIT_18 => X"100022012100102121082b40002108171216021502140213b5116b10b16c7100",
INIT_19 => X"ff2bf201002110003c012100102121082b21013e2b40002110f4212bf2010021",
INIT_1A => X"002110072184712156ac7100172a23505021002171740000002c71002b2c10f4",
INIT_1B => X"018c71000080015a00055fe0000021102188710021f4012171ff010521710056",
INIT_1C => X"736f6b6763383430343863676b6f7377006c0187002100e32a105090710021f1",
INIT_1D => X"702020200052206720200074202c0072626f202c000032200020616f432d0077",
INIT_1E => X"78206e007400676d6f006f002e6e726769006573640061742020006c20202000",
INIT_1F => X"00000000000000000000000000000000000020003a6874003a68740000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
